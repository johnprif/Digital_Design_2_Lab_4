library verilog;
use verilog.vl_types.all;
entity ADDER_8Bits_ADDSUB_vlg_vec_tst is
end ADDER_8Bits_ADDSUB_vlg_vec_tst;
