library verilog;
use verilog.vl_types.all;
entity Flag_Reg_vlg_vec_tst is
end Flag_Reg_vlg_vec_tst;
