library verilog;
use verilog.vl_types.all;
entity my_mux_2_1_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end my_mux_2_1_vlg_check_tst;
