library verilog;
use verilog.vl_types.all;
entity Flag_Reg_vlg_check_tst is
    port(
        FLAG_OUT        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Flag_Reg_vlg_check_tst;
