library verilog;
use verilog.vl_types.all;
entity my_mux_2_1_vlg_vec_tst is
end my_mux_2_1_vlg_vec_tst;
