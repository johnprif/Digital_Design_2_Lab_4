library verilog;
use verilog.vl_types.all;
entity REG_A_vlg_vec_tst is
end REG_A_vlg_vec_tst;
